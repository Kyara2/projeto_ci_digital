`timescale 1ns / 1ps

module button_interface_tb();

    // Sinais de entrada (reg) e sa�da (wire)
    reg clk;
    reg btn_in;
    wire btn_tick;

    // Instancia o m�dulo sob teste (UUT)
    button_interface uut (
        .clk(clk),
        .btn_in(btn_in),
        .btn_tick(btn_tick)
    );

    // Gera��o do Clock de 12 MHz
    // Per�odo: 1 / 12MHz = 83.33ns. Metade do ciclo = 41.66ns
    always begin
        #41.66 clk = ~clk;
    end

    initial begin
        // Inicializa��o
        clk = 0;
        btn_in = 1; // Bot�o solto (Active Low)
        
        $display("Iniciando simula��o...");
        #100;

        // --- Simula��o de Aperto de Bot�o com Ru�do (Bouncing) ---
        $display("Simulando ru�do de descida (bouncing)...");
        btn_in = 0; #100;
        btn_in = 1; #150;
        btn_in = 0; #200;
        btn_in = 1; #100;
        
        // Agora o bot�o estabiliza em 0 (pressionado)
        $display("Bot�o estabilizado em LOW. Aguardando tempo de debounce...");
        btn_in = 0;

        // Precisamos esperar mais de 1.200.000 ciclos. 
        // 1.200.000 * 83.33ns = ~100ms
        // Em simula��o, isso pode ser demorado. 
        // Se quiser testar r�pido, diminua o 'number_of_cycles' no c�digo original.
        #105000000; // Espera 105ms

        if (btn_tick) 
            $display("Sucesso: btn_tick detectado ap�s debounce!");
        else 
            $display("Erro: btn_tick n�o detectado.");

        #1000;

        // --- Simula��o de Soltura de Bot�o ---
        $display("Simulando soltura do bot�o...");
        btn_in = 1; 
        
        #105000000; // Espera mais 105ms para estabilizar em HIGH

        $display("Simula��o finalizada.");
        $finish;
    end

    // Opcional: Gerar arquivo para visualizar as ondas no GTKWave
    initial begin
        $dumpfile("button_interface_tb.vcd");
        $dumpvars(0, button_interface_tb);
    end

endmodule