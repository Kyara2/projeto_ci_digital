`timescale 1ns / 1ps


module ice_sugar (
	// input gpios  ------------
    input  wire clk,
	
	// buttons
    input  wire button_reset, 
    input  wire button_a,
	
	// receive uart
    input  wire rx,
	
	// output gpios ----------------
	// transmit uart
    output wire tx,
	
	// display with 4 digits
    output wire [6:0] seg,
    output wire [3:0] digits,
	
	// led rgb and external led
	output red, green, blue, test_button_led,
	
	// i2c interface
	inout wire i2c_scl,
	inout wire i2c_sda
);

	localparam DISPLAY_VALUE_BYTES = 2;
	
	localparam BYTES_FROM_DEBUG = 8; //15;
	localparam BYTES_TO_SEND_UART = BYTES_FROM_DEBUG*2 + 2;
	localparam BYTES_FROM_SENSOR = 2;

    wire button_reset_pressed;
    wire button_a_pressed;	
		
	wire [DISPLAY_VALUE_BYTES*8-1:0] display_value; 
	wire [15:0] rx_data;
	wire        rx_ready;
	wire [15:0] tx_data;
	
	wire tx_busy_total_signal;
	
	wire [BYTES_FROM_SENSOR*8-1:0] sensor_data;

	wire [BYTES_FROM_DEBUG*8-1:0] debug_bits;
    wire [(BYTES_FROM_DEBUG*2)*8-1:0] data_converted_to_ascii; // 4 nibbles convertidos para ASCII
	wire [BYTES_TO_SEND_UART*8-1:0] full_uart_frame; // 4 nibbles convertidos para ASCII
	wire [BYTES_TO_SEND_UART*8-1:0] frame_from_uart;
		
    assign debug_bits = 64'h01_23_45_67_89_AB_CD_EF; // for testing only
	//assign display_value = frame_from_uart[15:0];  // 16'h5678; // for testing only
	
	translate_hex_to_ascii #(.NUM_BYTES(BYTES_FROM_DEBUG)) converter (
		.data_in(debug_bits),
		.ascii_out(data_converted_to_ascii)
    );
	
	// Monta o frame: N caracteres de debug + \r\n(new line)
	assign full_uart_frame = {data_converted_to_ascii, 16'h0A0D};
	
	//assign display_value = sensor_data;  
	assign display_value = frame_from_uart[DISPLAY_VALUE_BYTES*8-1:0]; // for debug only
	
	// Se o mestre quer enviar 0, a FPGA puxa para 0. 
	// Se o mestre quer enviar 1, a FPGA solta (1'bz) e o resistor de 2.2k sobe a linha.
	// Se o mestre quer mandar 0, forçamos 0. Se quer mandar 1, soltamos (Z).
	// Se o mestre quer 0, a FPGA força 0. Se quer 1, a FPGA solta (1'bz).
	// Garante comportamento Open-Drain puro
	// Mude no topo ice_sugar.v:
	// Use buffers de dreno aberto explícitos
	//
	
	wire sda_in, sda_out, sda_dir;
	wire scl_in, scl_out, scl_dir;
	// Garante que o pino só vá para 0 ou Z (nunca force 1)
	
	
	//assign scl_dir = 1'b1; // button_a_pressed; //1'b1;
	//assign sda_dir = 1'b1; // button_a_pressed; // 1'b1;
	// Correção do Tri-state para I2C
	// Puxa para 0 apenas se a direção for saída (1) E o dado for 0.
	// Se o dado for 1 ou a direção for entrada (0), fica em Z.
	assign i2c_scl = (scl_dir && !scl_out) ? 1'b0 : 1'bz;
	assign i2c_sda = (sda_dir && !sda_out) ? 1'b0 : 1'bz;

	// As entradas continuam iguais
	assign scl_in = i2c_scl;
	assign sda_in = i2c_sda;
	

    // Instância para Reset (gera um pulso de reset)
    button_interface btn_reset (
        .clk(clk),
        .btn_in(button_reset),
        .btn_tick(button_reset_pressed)
    );

    // Instância para Send (gera um pulso para enviar)
    button_interface btn_a (
        .clk(clk),
        .btn_in(button_a),
        .btn_tick(button_a_pressed)
    );
	
	// leds
	leds_interface leds (
		.clk(clk),
		.reset(button_reset_pressed),
		.signal(button_a_pressed),
		.red(red),
		.green(green),
		.blue(blue),
		.test_led(test_button_led)
	);
	
	display_four_digits display_inst (
			.clk(clk),
			.reset(button_reset_pressed),
			.start_signal(button_a_pressed),
			//.start_signal(1'b1),
			//.input_value(display_value), // Mostra os 2 bytes acumulados
			.input_value(display_value),
			.seg(seg),
			.digits(digits)
		);
	
	
	uart_controller #(.BYTES(BYTES_TO_SEND_UART)) uart_controller_main (
        .clk(clk),
        .reset_n(!button_reset_pressed),
        //.data_to_send(input_data),
		.data_to_send(full_uart_frame),
        .start_tx(button_a_pressed),
		//.start_tx(1'b1),
        .data_received(frame_from_uart),
        .rx_done_tick(rx_ready),
        .tx_busy_total(tx_busy_total_signal),
        .rx(rx),
        .tx(tx)
    );
    
	
	
	
	// Instancia o seu controlador que gerencia o Master e o Sensor
	
	i2c_controller #(
		.BYTES_FROM_DATA(BYTES_FROM_SENSOR),
		.BYTES_FROM_DEBUG(BYTES_FROM_DEBUG)
	) user_app (
		.clk(clk),
		.reset(button_reset_pressed), 
		.start_pulse(button_a_pressed), 
		.sda_in(sda_in), .scl_in(scl_in),
		.sda_out(sda_out), .scl_out(scl_out),
		.sda_dir(sda_dir), .scl_dir(scl_dir),
		//.debug_bits(debug_bits),
		.sensor_data(sensor_data)
	);
	
	
	wire [31:0] x1, x2, x3, pc_out, instr_out, alu_out, reg_wirte_out;
	
	cpu_top RV32I (
		.clk(clk),
		.reset(button_reset_pressed),
		.x1(x1),
		.x2(x2),
		.x3(x3),
		.pc_out(pc_out),
		.instr_out(instr_out),
		.alu_out(alu_out),
		.reg_write_out(reg_write_out)
	);
endmodule




